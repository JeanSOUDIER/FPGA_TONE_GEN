library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
	generic(constant ROM_SIZE_X : natural := 5; constant ROM_SIZE_Y : natural := 2; constant DATA_WIDTH : natural := 32);
	port (
		CLK, RST : std_logic;
		ADDR : in std_logic_vector((ROM_SIZE_X)*(ROM_SIZE_Y)-1 downto 0);
		Q : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity;

architecture bhv of ROM is
type rom_type is array (0 to 2**((ROM_SIZE_X)*(ROM_SIZE_Y))-1) of integer;
constant data : rom_type :=(
--Sine
0	,
52701887	,
105372029	,
157978698	,
210490206	,
262874924	,
315101295	,
367137861	,
418953277	,
470516331	,
521795963	,
572761286	,
623381598	,
673626408	,
723465452	,
772868706	,
821806413	,
870249095	,
918167572	,
965532978	,
1012316784	,
1058490808	,
1104027237	,
1148898640	,
1193077991	,
1236538675	,
1279254515	,
1321199780	,
1362349204	,
1402677999	,
1442161874	,
1480777044	,
1518500250	,
1555308768	,
1591180425	,
1626093616	,
1660027308	,
1692961062	,
1724875040	,
1755750017	,
1785567396	,
1814309216	,
1841958164	,
1868497585	,
1893911494	,
1918184580	,
1941302225	,
1963250501	,
1984016188	,
2003586779	,
2021950483	,
2039096241	,
2055013723	,
2069693341	,
2083126254	,
2095304369	,
2106220351	,
2115867625	,
2124240380	,
2131333571	,
2137142927	,
2141664948	,
2144896909	,
2146836866	,
2147483647	,
2146836866	,
2144896909	,
2141664948	,
2137142927	,
2131333571	,
2124240380	,
2115867625	,
2106220351	,
2095304369	,
2083126254	,
2069693341	,
2055013723	,
2039096241	,
2021950483	,
2003586779	,
1984016188	,
1963250501	,
1941302225	,
1918184580	,
1893911494	,
1868497585	,
1841958164	,
1814309216	,
1785567396	,
1755750017	,
1724875040	,
1692961062	,
1660027308	,
1626093616	,
1591180425	,
1555308768	,
1518500250	,
1480777044	,
1442161874	,
1402677999	,
1362349204	,
1321199780	,
1279254515	,
1236538675	,
1193077991	,
1148898640	,
1104027237	,
1058490808	,
1012316784	,
965532978	,
918167572	,
870249095	,
821806413	,
772868706	,
723465452	,
673626408	,
623381598	,
572761286	,
521795963	,
470516331	,
418953277	,
367137861	,
315101295	,
262874924	,
210490206	,
157978698	,
105372029	,
52701887	,
1	,
-52701887	,
-105372029	,
-157978698	,
-210490206	,
-262874924	,
-315101295	,
-367137861	,
-418953277	,
-470516331	,
-521795963	,
-572761286	,
-623381598	,
-673626408	,
-723465452	,
-772868706	,
-821806413	,
-870249095	,
-918167572	,
-965532978	,
-1012316784	,
-1058490808	,
-1104027237	,
-1148898640	,
-1193077991	,
-1236538675	,
-1279254515	,
-1321199780	,
-1362349204	,
-1402677999	,
-1442161874	,
-1480777044	,
-1518500250	,
-1555308768	,
-1591180425	,
-1626093616	,
-1660027308	,
-1692961062	,
-1724875040	,
-1755750017	,
-1785567396	,
-1814309216	,
-1841958164	,
-1868497585	,
-1893911494	,
-1918184580	,
-1941302225	,
-1963250501	,
-1984016188	,
-2003586779	,
-2021950483	,
-2039096241	,
-2055013723	,
-2069693341	,
-2083126254	,
-2095304369	,
-2106220351	,
-2115867625	,
-2124240380	,
-2131333571	,
-2137142927	,
-2141664948	,
-2144896909	,
-2146836866	,
-2147483647	,
-2146836866	,
-2144896909	,
-2141664948	,
-2137142927	,
-2131333571	,
-2124240380	,
-2115867625	,
-2106220351	,
-2095304369	,
-2083126254	,
-2069693341	,
-2055013723	,
-2039096241	,
-2021950483	,
-2003586779	,
-1984016188	,
-1963250501	,
-1941302225	,
-1918184580	,
-1893911494	,
-1868497585	,
-1841958164	,
-1814309216	,
-1785567396	,
-1755750017	,
-1724875040	,
-1692961062	,
-1660027308	,
-1626093616	,
-1591180425	,
-1555308768	,
-1518500250	,
-1480777044	,
-1442161874	,
-1402677999	,
-1362349204	,
-1321199780	,
-1279254515	,
-1236538675	,
-1193077991	,
-1148898640	,
-1104027237	,
-1058490808	,
-1012316784	,
-965532978	,
-918167572	,
-870249095	,
-821806413	,
-772868706	,
-723465452	,
-673626408	,
-623381598	,
-572761286	,
-521795963	,
-470516331	,
-418953277	,
-367137861	,
-315101295	,
-262874924	,
-210490206	,
-157978698	,
-105372029	,
-52701887	,
--Square
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
-2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
2147483647	,
--Triangle
-2147483647	,
-2113929216	,
-2080374784	,
-2046820352	,
-2013265920	,
-1979711488	,
-1946157056	,
-1912602624	,
-1879048192	,
-1845493760	,
-1811939328	,
-1778384896	,
-1744830464	,
-1711276032	,
-1677721600	,
-1644167168	,
-1610612736	,
-1577058304	,
-1543503872	,
-1509949440	,
-1476395008	,
-1442840576	,
-1409286144	,
-1375731712	,
-1342177280	,
-1308622848	,
-1275068416	,
-1241513984	,
-1207959552	,
-1174405120	,
-1140850688	,
-1107296256	,
-1073741824	,
-1040187392	,
-1006632960	,
-973078528	,
-939524096	,
-905969664	,
-872415232	,
-838860800	,
-805306368	,
-771751936	,
-738197504	,
-704643072	,
-671088640	,
-637534208	,
-603979776	,
-570425344	,
-536870912	,
-503316480	,
-469762048	,
-436207616	,
-402653184	,
-369098752	,
-335544320	,
-301989888	,
-268435456	,
-234881024	,
-201326592	,
-167772160	,
-134217728	,
-100663296	,
-67108864	,
-33554432	,
0	,
33554432	,
67108864	,
100663296	,
134217728	,
167772160	,
201326592	,
234881024	,
268435456	,
301989888	,
335544320	,
369098752	,
402653184	,
436207616	,
469762048	,
503316480	,
536870912	,
570425344	,
603979776	,
637534208	,
671088640	,
704643072	,
738197504	,
771751936	,
805306368	,
838860800	,
872415232	,
905969664	,
939524096	,
973078528	,
1006632960	,
1040187392	,
1073741824	,
1107296256	,
1140850688	,
1174405120	,
1207959552	,
1241513984	,
1275068416	,
1308622848	,
1342177280	,
1375731712	,
1409286144	,
1442840576	,
1476395008	,
1509949440	,
1543503872	,
1577058304	,
1610612736	,
1644167168	,
1677721600	,
1711276032	,
1744830464	,
1778384896	,
1811939328	,
1845493760	,
1879048192	,
1912602624	,
1946157056	,
1979711488	,
2013265920	,
2046820352	,
2080374784	,
2113929216	,
2147483647	,
2113929216	,
2080374784	,
2046820352	,
2013265920	,
1979711488	,
1946157056	,
1912602624	,
1879048192	,
1845493760	,
1811939328	,
1778384896	,
1744830464	,
1711276032	,
1677721600	,
1644167168	,
1610612736	,
1577058304	,
1543503872	,
1509949440	,
1476395008	,
1442840576	,
1409286144	,
1375731712	,
1342177280	,
1308622848	,
1275068416	,
1241513984	,
1207959552	,
1174405120	,
1140850688	,
1107296256	,
1073741824	,
1040187392	,
1006632960	,
973078528	,
939524096	,
905969664	,
872415232	,
838860800	,
805306368	,
771751936	,
738197504	,
704643072	,
671088640	,
637534208	,
603979776	,
570425344	,
536870912	,
503316480	,
469762048	,
436207616	,
402653184	,
369098752	,
335544320	,
301989888	,
268435456	,
234881024	,
201326592	,
167772160	,
134217728	,
100663296	,
67108864	,
33554432	,
0	,
-33554432	,
-67108864	,
-100663296	,
-134217728	,
-167772160	,
-201326592	,
-234881024	,
-268435456	,
-301989888	,
-335544320	,
-369098752	,
-402653184	,
-436207616	,
-469762048	,
-503316480	,
-536870912	,
-570425344	,
-603979776	,
-637534208	,
-671088640	,
-704643072	,
-738197504	,
-771751936	,
-805306368	,
-838860800	,
-872415232	,
-905969664	,
-939524096	,
-973078528	,
-1006632960	,
-1040187392	,
-1073741824	,
-1107296256	,
-1140850688	,
-1174405120	,
-1207959552	,
-1241513984	,
-1275068416	,
-1308622848	,
-1342177280	,
-1375731712	,
-1409286144	,
-1442840576	,
-1476395008	,
-1509949440	,
-1543503872	,
-1577058304	,
-1610612736	,
-1644167168	,
-1677721600	,
-1711276032	,
-1744830464	,
-1778384896	,
-1811939328	,
-1845493760	,
-1879048192	,
-1912602624	,
-1946157056	,
-1979711488	,
-2013265920	,
-2046820352	,
-2080374784	,
-2113929216	,
--Rampe
-2147483647	,
-2130706432	,
-2113929216	,
-2097152000	,
-2080374784	,
-2063597568	,
-2046820352	,
-2030043136	,
-2013265920	,
-1996488704	,
-1979711488	,
-1962934272	,
-1946157056	,
-1929379840	,
-1912602624	,
-1895825408	,
-1879048192	,
-1862270976	,
-1845493760	,
-1828716544	,
-1811939328	,
-1795162112	,
-1778384896	,
-1761607680	,
-1744830464	,
-1728053248	,
-1711276032	,
-1694498816	,
-1677721600	,
-1660944384	,
-1644167168	,
-1627389952	,
-1610612736	,
-1593835520	,
-1577058304	,
-1560281088	,
-1543503872	,
-1526726656	,
-1509949440	,
-1493172224	,
-1476395008	,
-1459617792	,
-1442840576	,
-1426063360	,
-1409286144	,
-1392508928	,
-1375731712	,
-1358954496	,
-1342177280	,
-1325400064	,
-1308622848	,
-1291845632	,
-1275068416	,
-1258291200	,
-1241513984	,
-1224736768	,
-1207959552	,
-1191182336	,
-1174405120	,
-1157627904	,
-1140850688	,
-1124073472	,
-1107296256	,
-1090519040	,
-1073741824	,
-1056964608	,
-1040187392	,
-1023410176	,
-1006632960	,
-989855744	,
-973078528	,
-956301312	,
-939524096	,
-922746880	,
-905969664	,
-889192448	,
-872415232	,
-855638016	,
-838860800	,
-822083584	,
-805306368	,
-788529152	,
-771751936	,
-754974720	,
-738197504	,
-721420288	,
-704643072	,
-687865856	,
-671088640	,
-654311424	,
-637534208	,
-620756992	,
-603979776	,
-587202560	,
-570425344	,
-553648128	,
-536870912	,
-520093696	,
-503316480	,
-486539264	,
-469762048	,
-452984832	,
-436207616	,
-419430400	,
-402653184	,
-385875968	,
-369098752	,
-352321536	,
-335544320	,
-318767104	,
-301989888	,
-285212672	,
-268435456	,
-251658240	,
-234881024	,
-218103808	,
-201326592	,
-184549376	,
-167772160	,
-150994944	,
-134217728	,
-117440512	,
-100663296	,
-83886080	,
-67108864	,
-50331648	,
-33554432	,
-16777216	,
0	,
16777216	,
33554432	,
50331648	,
67108864	,
83886080	,
100663296	,
117440512	,
134217728	,
150994944	,
167772160	,
184549376	,
201326592	,
218103808	,
234881024	,
251658240	,
268435456	,
285212672	,
301989888	,
318767104	,
335544320	,
352321536	,
369098752	,
385875968	,
402653184	,
419430400	,
436207616	,
452984832	,
469762048	,
486539264	,
503316480	,
520093696	,
536870912	,
553648128	,
570425344	,
587202560	,
603979776	,
620756992	,
637534208	,
654311424	,
671088640	,
687865856	,
704643072	,
721420288	,
738197504	,
754974720	,
771751936	,
788529152	,
805306368	,
822083584	,
838860800	,
855638016	,
872415232	,
889192448	,
905969664	,
922746880	,
939524096	,
956301312	,
973078528	,
989855744	,
1006632960	,
1023410176	,
1040187392	,
1056964608	,
1073741824	,
1090519040	,
1107296256	,
1124073472	,
1140850688	,
1157627904	,
1174405120	,
1191182336	,
1207959552	,
1224736768	,
1241513984	,
1258291200	,
1275068416	,
1291845632	,
1308622848	,
1325400064	,
1342177280	,
1358954496	,
1375731712	,
1392508928	,
1409286144	,
1426063360	,
1442840576	,
1459617792	,
1476395008	,
1493172224	,
1509949440	,
1526726656	,
1543503872	,
1560281088	,
1577058304	,
1593835520	,
1610612736	,
1627389952	,
1644167168	,
1660944384	,
1677721600	,
1694498816	,
1711276032	,
1728053248	,
1744830464	,
1761607680	,
1778384896	,
1795162112	,
1811939328	,
1828716544	,
1845493760	,
1862270976	,
1879048192	,
1895825408	,
1912602624	,
1929379840	,
1946157056	,
1962934272	,
1979711488	,
1996488704	,
2013265920	,
2030043136	,
2046820352	,
2063597568	,
2080374784	,
2097152000	,
2113929216	,
2130706432	
);
begin
	process(CLK, RST)
	begin
		if (RST = '0') then
			Q <= (others=>'0');
		elsif (rising_edge(CLK)) then
			Q <= std_logic_vector(to_signed(data(to_integer(unsigned(ADDR))),DATA_WIDTH));
		end if;
	end process;
end architecture;
